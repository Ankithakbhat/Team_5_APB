`include "apb_test.sv"