interface apb_intrf(bit clk, bit rst);




endinterface