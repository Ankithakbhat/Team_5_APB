`include "base_test.sv"
`include "read_error.sv"
`include "write_error.sv"
`include "write.sv"
`include "read.sv"
`include "write_read_0.sv"
`include "write_read_1.sv"
`include "alternate_read_write.sv"
