`include "apb_sequence_item.sv"
