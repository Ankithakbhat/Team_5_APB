`define AW 5
`define DW 32
`define SW 4